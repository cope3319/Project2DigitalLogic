module segToDec(seg1,seg2,dig1,dig2)
input [7:0] seg1;
input [7:0] seg2;
output [3:0] dig1;
output [3:0] dig2;

always @*
begin
    casex(seg1[7:0])
        8'b11000000 : dig1 = 4'b0000; //0
        8'b11111001 : dig1 = 4'b0001; //1
        8'b10100100 : dig1 = 4'b0010; //2
        8'b10110000 : dig1 = 4'b0011; //3
        8'b10011001 : dig1 = 4'b0100; //4
        8'b10010010 : dig1 = 4'b0101; //5
        8'b10000010 : dig1 = 4'b0110; //6
        8'b11111000 : dig1 = 4'b0111; //7
        8'b10000000 : dig1 = 4'b1000; //8
        8'b10010000 : dig1 = 4'b1001; //9
    endcase
    casex(seg2[7:0])
        8'b11000000 : dig2 = 4'b0000; //0
        8'b11111001 : dig2 = 4'b0001; //1
        8'b10100100 : dig2 = 4'b0010; //2
        8'b10110000 : dig2 = 4'b0011; //3
        8'b10011001 : dig2 = 4'b0100; //4
        8'b10010010 : dig2 = 4'b0101; //5
        8'b10000010 : dig2 = 4'b0110; //6
        8'b11111000 : dig2 = 4'b0111; //7
        8'b10000000 : dig2 = 4'b1000; //8
        8'b10010000 : dig2 = 4'b1001; //9
    endcase
end
end