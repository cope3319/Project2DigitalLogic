module monthDayCalc(data,month,day)


endmodule